module TTT()

  
endmodule
