module TTT()
hihi
