module game(clk, key_data, IsItMain, board, IsItRight)
  input clk;
  input key_data;
  input IsItMain;
  
