module TTT()

  
endmodule