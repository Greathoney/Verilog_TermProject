module source(CLOCK, RESET)

endmodule

