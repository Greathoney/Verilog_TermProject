module
sdfsd
