module TTT()



//input 
