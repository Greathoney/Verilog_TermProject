module TTT(CLOCK, RESET)

endmodule
