module TTT()
